library IEEE;

use IEEE.std_logic_1164.all;

use IEEE.numeric_std.all;

-- We are programming on VHDL. This is a VHDL file.

entity multiplicator is
  port(
    instruction_i : in  std_logic_vector(31 downto 0);
    rs1_i         : in  std_logic_vector(31 downto 0);
    rs2_i         : in  std_logic_vector(31 downto 0);
    result_o      : out std_logic_vector(31 downto 0);
    icc_o         : out std_logic_vector(3 downto 0)
    );
end;



architecture multiplicator_arq of multiplicator is
  constant UMUL_OPCODE : std_logic_vector(5 downto 0) := "011010";
  constant SMUL_OPCODE : std_logic_vector(5 downto 0) := "011011";

  signal operand2 : std_logic_vector(31 downto 0) := (others => '0');
  signal result   : std_logic_vector(31 downto 0) := (others => '0');


  function debug_vector_as_string (a : std_logic_vector) return string is
    variable b    : string (1 to a'length) := (others => NUL);
    variable stri : integer                := 1;
  begin
    for i in a'range loop
      b(stri) := std_logic'image(a((i)))(2);
      stri    := stri+1;
    end loop;
    return b;
  end function;

  function signed_multiplication(L, R : std_logic_vector(31 downto 0)) return std_logic_vector is
    variable ret : std_logic_vector(63 downto 0);
  begin
    ret := std_logic_vector(signed(L) * signed(R));
    return ret(31 downto 0);
  end;


  function unsigned_multiplication(L, R : std_logic_vector(31 downto 0)) return std_logic_vector is
    variable ret : std_logic_vector(63 downto 0);
  begin
    ret := std_logic_vector(unsigned(L) * unsigned(R));
    return ret(31 downto 0);
  end;


begin
  -- operand2 := if (i = 0) then r[rs2] else sign_extend(simm13); INFO: (A)
  --
  -- INFO: (B)
  -- if (UMUL or UMULcc) then
  --   (Y, result) ← multiply_unsigned(r[rs1], operand2);
  -- else if (SMUL or SMULcc) then
  --   (Y, result) ← multiply_signed(r[rs1], operand2);
  --
  -- next;
  --
  -- if (rd ≠ 0) then INFO: We assume always TRUE
  --   r[rd] ← result; INFO: (C)
  --
  -- if (UMULcc or SMULcc) then ( INFO: Always TRUE
  --   N ← result<31>; INFO: (D)
  --
  --   Z ← if (result = 0) then 1 else 0; INFO: (E)
  --
  --   INFO: (F)
  --   V ← 0;
  --
  --   INFO: (G)
  --   C ← 0
  -- );

  -- BEGIN: (A)
  -- Check the 13bit of `instruction_i`
  process(instruction_i, rs1_i, rs2_i)
  begin
    if instruction_i(13) = '0' then
      operand2 <= rs2_i;
    else
      -- Move the last 13bits of `instruction_i` to `operand2`
      operand2 <= (31 downto 13 => '0') & instruction_i(12 downto 0);
    end if;
  end process;

  -- BEGIN: (B)
  -- Calculate the multiplication and assing to `result`
  result <= signed_multiplication(rs1_i, operand2) when (instruction_i(24 downto 19) = SMUL_OPCODE) else
            unsigned_multiplication(rs1_i, operand2) when (instruction_i(24 downto 19) = UMUL_OPCODE) else
            (others => '0');  -- In reality this should never happen...

  -- BEGIN: (C)
  -- Assing the result to `result_o`
  result_o <= result;

  -- BEGIN: (D)
  -- Assing the 31bit of `result` to `icc_o(3)`
  icc_o(3) <= result(31);

  -- BEGIN: (E)
  -- Assing the 0 or 1 to `icc_o`
  icc_o(2) <= '1' when result = "00000000000000000000000000000000" else '0';

  -- BEGIN: (F)
  -- Assing the V to `icc_o`
  -- process(rs1_i, operand2, result)
  -- begin
  --   report "RS1:      " & debug_vector_as_string(rs1_i);
  --   report "operand2: " & debug_vector_as_string(operand2);
  --   report "result:   " & debug_vector_as_string(result);
  --   report "-----------";
  -- end process;

  icc_o(1) <= '0';

  -- BEGIN: (G)
  -- Assing the C to `icc_o`
  icc_o(0) <= '0';

end;
